Colpitts Oscillator
*
* @brief : Colpitts Oscillator 
* @author : S.Dusausay
*

*.subckt COLPITTS C E 
.include ./2N2222.cir

* Av
VCC A 0 DC=15
RB2 A B 150k
RB1 B 0 22k
Cde B 0 100n
Q1  C B E 2N2222
RE  E 0 1040

* b(w)
L1  A C 220n
C1  C E 30p
C2  E 0 30p 

*.ends

.control
tran 10p 0.5u 0u 10p
plot V(E) V(C)
.endc
.end
