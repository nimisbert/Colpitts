
.model 2N2222 NPN( 
+ IS=1E-14 
+ VAF=100 
+ BF=200 
+ IKF=0.3 
+ XTB=1.5 
+ BR=3 
+ CJC=8E-12 
+ CJE=25E-12 
+ TR=100E-9 
+ TF=400E-12 
+ ITF=1 
+ VTF=2 
+ XTF=3 
+ RB=10 
+ RC=.3 
+ RE=.2) 
*+ Vceo=30 
*+ Icrating=800m 
*+ mfg=Philips)
